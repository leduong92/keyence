[HD]
CPDF_B  V1.3
LINK    1
FILE  0
DEF_CNT  0
REF_CNT  0
[FILE]
[CLASS]
[MEMBER]
[OBJECT]
[CONST]
